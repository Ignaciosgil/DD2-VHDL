library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity master_spi_4_hilos is
port(nRst:     in     std_logic;
     clk:      in     std_logic;                       -- 50 MHz   (IMPORTANTE)
     -- Ctrl_SPI
     start:    in     std_logic;                       -- Orden de ejecucion (si rdy = 1 ) => rdy  <= 0 hasta fin, cuando rdy <= 1
     nWR_RD:   in     std_logic;                       -- Escritura (0) o lectura (1)
     dir_reg:  in     std_logic_vector(6 downto 0);    -- direccion de acceso; si bit 7 a 1 (autoincremento) y RD, se considera el valor de long
     dato_wr:  in     std_logic_vector(7 downto 0);    -- dato a escribir (solo escrituras de 1 bit
     dato_rd:  buffer std_logic_vector(7 downto 0);    -- valor del byte leido
     ena_rd:   buffer std_logic;                       -- valida a nivel alto a dato_rd -> Ignorar en operacion de escritura
     rdy:      buffer std_logic;                       -- unidad preparada para aceptar start
     -- bus SPI
     nCS:      buffer std_logic;                      -- chip select
     SPC:      buffer std_logic;                      -- clock SPI
     SDI:      in     std_logic;                      -- Master Data input (connected to slave SDO)
     SDO:      buffer std_logic);                     -- Master Data Output (connected to slave SDI)         NO hay que sincronizar la se�al, p
     
end entity;

architecture rtl of master_spi_4_hilos is
 --Reloj del bus
 signal cnt_SPC:     std_logic_vector(2 downto 0);
 signal fdc_cnt_SPC: std_logic;
 signal SPC_posedge: std_logic;
 signal SPC_negedge: std_logic;

 constant SPC_LH: natural := 5; 
 
 -- Contador de bits y bytes transmitidos
 signal cnt_bits_SPC: std_logic_vector(5 downto 0);

 -- Sincro SDI y Registro de transmision y recepcion
 signal SDI_meta, SDI_syn: std_logic;
 signal reg_SPI: std_logic_vector(16 downto 0);

 -- Para el control
 signal no_bytes: std_logic_vector(2 downto 0); 
 signal fin: std_logic;

begin
  -- Generacion de nCS:
  process(nRst, clk)
  begin
    if nRst = '0' then
      nCS <= '1';

    elsif clk'event and clk = '1' then
      if start = '1' and nCS = '1' then
        nCS <= '0';

      elsif fin = '1' then
        nCS <= '1';

      end if;
    end if;
  end process;
  
  rdy <= nCS;

  -- Generacion de SPC: FLIP FLOP TIPO T
  -- SPC se�al registrada
  process(nRst, clk)
  begin
    if nRst = '0' then
      cnt_SPC <= (0 => '1', others => '0');   -- Porque comienza desde 10  -> 2 decimal
      SPC <= '1';

    elsif clk'event and clk = '1' then
      if nCS = '1' then 
        cnt_SPC <= (0 => '1', others => '0');
        SPC <= '1';

      elsif fdc_cnt_SPC = '1' then   -- cuando el contador cnt_SPC llegue a 5 cambia el nivel de la se�al  (periodo del reloj = 10 cnt_SPC)
        SPC <= not SPC;
        cnt_SPC <= (0 => '1', others => '0');  -- Y aqui comienza desde 1

      else
        cnt_SPC <= cnt_SPC + 1;

      end if;
    end if;
  end process;

  --Esto hace que el reloj sea cuadrado =t a NA y a NB
  fdc_cnt_SPC <= '1' when cnt_SPC = SPC_LH else           -- cada 100 ns
                 '0';

  --Flanco de subida y flanco de bajada 

  SPC_posedge <= SPC when cnt_SPC = 1 else       -- Cuando el estado de cuenta vale 1, SPC siempre vale 1
                 '0'; 

  SPC_negedge <= not SPC when cnt_SPC = 1 else   -- Siempre valdra cero
                 '0'; 

  -- Cuenta bits y bytes:
  process(nRst, clk)
  begin
    if nRst = '0' then
      cnt_bits_SPC <= (others => '0');
      
    elsif clk'event and clk = '1' then  
      if SPC_posedge = '1' then			--SPC cuenta bits en los flancos de subida 
        cnt_bits_SPC <= cnt_bits_SPC + 1;

      elsif nCS = '1' then               -- Se resetea cuando termina la transferencia nCs = '1'
        cnt_bits_SPCcnt_bits_SPC <= (others => '0');

      end if;
    end if;
  end process;

  -- Registro
  process(nRst, clk)
  begin
    if nRst = '0' then
      reg_SPI <= (others => '0');
      SDI_syn <= '0';
      SDI_meta <= '0';

    elsif clk'event and clk = '1' then  
      SDI_meta <= SDI;					-- Es el bus que usa el master para enviar datos al esclavo
      SDI_syn <= SDI_meta;				-- Estoy sincronizando la se�al,asi evito los glitches
      
      if start = '1' and nCS = '1' then  		-- Empiezo una transferencia 
        reg_SPI <= '0'& nWR_RD & dir_reg & dato_wr;  	-- Guardo si es lectura/escritura, la dir del reg donde opero, y el dato (si se trata de una escritura)
 
      elsif SPC_negedge = '1' then 			-- El master lee lo que le manda el esclavo
        reg_SPI(16 downto 1) <= reg_SPI(15 downto 0);   -- Guardo los 2 bytes de lectura en la parte mas alta del registro

      elsif SPC_posedge = '1' then			-- El master escribe en el bit de menos peso   ???
        reg_SPI(0) <= SDI_syn;

      end if;
    end if;
  end process;

--Habilitacion de lectura 
  ena_rd <= (not nCS and fin) when cnt_bits_SPC(5 downto 3) =  no_bytes else  --COMPLETAR
            SPC_negedge       when cnt_bits_SPC(5 downto 3) > 1  and cnt_bits_SPC(2 downto 0) = 7 else  --COMPLETAR  El byte esta completo
            '0';

  dato_rd <= reg_SPI(7 downto 0);	--valor del dato leido 

  SDO <= reg_SPI(16);	--voy mostrando el bit mas significativo

  -- Control heuristico
  process(nRst, clk)
  begin
    if nRst = '0' then
      no_bytes <= (others => '0');

    elsif clk'event and clk = '1' then  
      if start = '1' and nCS = '1' then
        if nWR_RD = '0' then		--indica si es lectura o escritura, si es 0 es una escritura el no_bytes que voy a escribir es 
          no_bytes <= "010" ;           -- si se trata de una escritura tengo 1 byte con la dir reg y 1 byte con los datos

        else
          no_bytes <= "011" ;          -- si se trata de una lectura tengo 1 byte con la dir reg y 2 bytes con los datos que se van a leer

        end if;
      end if;
    end if;
  end process;

  ---Se va si me encuentro en una escritura se realicen 2 bytes y si me encuentro en una lectura se realicen 3 bytes   ???? no seria escritura uno lectura dos
  fin <= '1' when cnt_bits_SPC(5 downto 3) = no_bytes else 
         '0';
 
end rtl;
